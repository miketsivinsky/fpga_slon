//------------------------------------------------------------------------------
//	Project:       slon03
//	Description:   The Second Xilinx slonick (slon02 - is a Pin Planning Project)
//------------------------------------------------------------------------------

`ifndef SLON_03_SVH
`define SLON_03_SVH


//******************************************************************************
//******************************************************************************
package slon03_lib;

//------------------------------------------------------------------------------
//    Settings
//

parameter integer GREEN_LED_NUM = 4;

endpackage : slon03_lib


`endif // SLON_03_SVH

