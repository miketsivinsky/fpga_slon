//------------------------------------------------------------------------------
//	Project:       slon01
//	Description:   The First Xilinx slonick
//------------------------------------------------------------------------------

//******************************************************************************
//******************************************************************************
module slon01
(
    output bit [7:4] ledGreen
);

//------------------------------------------------------------------------------
//    Settings
//

//------------------------------------------------------------------------------
//    Types
//

//------------------------------------------------------------------------------
//    Objects
//

//------------------------------------------------------------------------------
//    Functions and Tasks
//

//------------------------------------------------------------------------------
//     Logic
//

assign ledGreen = 4'b1010;

endmodule : slon01